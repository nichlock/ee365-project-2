library ieee;
use ieee.std_logic_1164.all;

package values is
	constant N: integer :=6;	-- must not be more than 6 for the DE0_Nano board			 
end package values;